
module Lab1_sys (
	clk_clk,
	pio_0_external_connection_export,
	reset_reset_n,
	pio_1_external_connection_export);	

	input		clk_clk;
	output	[7:0]	pio_0_external_connection_export;
	input		reset_reset_n;
	input		pio_1_external_connection_export;
endmodule
