
module Lab1_sys (
	clk_clk,
	pio_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output		pio_0_external_connection_export;
	input		reset_reset_n;
endmodule
